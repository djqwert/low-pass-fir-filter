library ieee;
use ieee.std_logic_1164.all;

entity reg is 
	generic(N: natural := 16);
	port(
		d: in std_logic_vector(N-1 downto 0);
		q: out std_logic_vector(N-1 downto 0);
		clk: in std_logic;
		rst: in std_logic;
		en: in std_logic
	);
end reg;

architecture bhv of reg is
begin

	
	process(clk,rst) 
	begin
		if rst = '0' then
			q <= (others => '0');
		elsif rising_edge(clk) then
			if en = '1' then
				q <= d;
			end if;
		end if;
	end process;

end bhv;